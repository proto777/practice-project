module inverter(in, out);

input in;
output out;

assign in = ~out ;

endmodule